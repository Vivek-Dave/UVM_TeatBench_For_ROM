
`include "interface.sv"
`include "tb_pkg.sv"
module top;
  import uvm_pkg::*;
  import tb_pkg::*;
  
  bit clk; // external signal declaration
  //----------------------------------------------------------------------------
  intf i_intf(clk);
  //----------------------------------------------------------------------------

  //----------------------------------------------------------------------------
  ROM DUT(.addr(i_intf.addr),
          .rd  (i_intf.rd),
          .out (i_intf.out),
          .clk (i_intf.clk),
          .rst(i_intf.rst)
         );
  //----------------------------------------------------------------------------               
  
  initial begin
    clk<=0;
  end

  always #5 clk=~clk;
  
  //----------------------------------------------------------------------------
  initial begin
    $dumpfile("dumpfile.vcd");
    $dumpvars;
  end
  //----------------------------------------------------------------------------

  //----------------------------------------------------------------------------
  initial begin
    uvm_config_db#(virtual intf)::set(uvm_root::get(),"","vif",i_intf);
  end
  //----------------------------------------------------------------------------

  //----------------------------------------------------------------------------
  initial begin
    run_test("rom_test");
  end
  //----------------------------------------------------------------------------
endmodule

