
`ifndef TB_PKG
`define TB_PKG
`include "uvm_macros.svh"
package tb_pkg;
 import uvm_pkg::*;
 `include "rom_sequence_item.sv"        // transaction class
 `include "rom_sequence.sv"             // sequence class
 `include "rom_sequencer.sv"            // sequencer class
 `include "rom_driver.sv"               // driver class
 `include "rom_monitor.sv"
 `include "rom_agent.sv"                // agent class  
 `include "rom_coverage.sv"             // coverage class
 `include "rom_scoreboard.sv"           // scoreboard class
 `include "rom_env.sv"                  // environment class

 `include "rom_test.sv"                 // test
endpackage
`endif 


